`ifndef __AXI_TYPEDEF_SVH__
`define	__AXI_TYPEDEF_SVH__

`define AXI_ADDR_WIDTH	64
`define AXI_DATA_WIDTH	32
`define AXI_ID_WIDTH	16
`define INDEX_WIDTH	4

`endif
