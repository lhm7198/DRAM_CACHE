`ifndef __FIFO_TYPEDEF_SVH__
`define	__FIFO_TYPEDEF_SVH__

`define FIFO_DATA_WIDTH		8
`define FIFO_HEIGHT		8
`define FIFO_A_FULL_THRH	6
`define FIFO_A_EMPTY_THR	2

`endif
